module and_gate(input logic [31:0] a, b, 
					output logic [31:0] c);

	assign c = a & b;

endmodule